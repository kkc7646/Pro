library ieee;
use ieee.std_logic_1164.all;
use IEEE.NUMERIC_STD.ALL;

entity memory is
	port(A			                  : in  std_logic_vector(15 downto 0);
			 Din                      : in std_logic_vector(15 downto 0);		
			 clock,mem_Write,mem_read : in  std_logic;
			 Dout				              : out std_logic_vector(15 downto 0));
end memory;

architecture Structure of memory is
type memory_16 is array (65535 downto 0) of std_logic_vector (15 downto 0);------------1kB of memory
signal T:memory_16 :=(0 => "1000001000000001",  ---JAL R1 0001H
											1 => "0100100110000101",  ---LW  R4 R6 0005H
											2 => "0001110000111101",  ---ADI R6 R0 111101B
											3 => "0100110110000101",  ---LW
											4 => "0100001101010101",  ---LW
											5 => "0001000010000000",  ---ADI
											6 => "0010000001011000",  ---NDU
											7 => "0010011011011000",  ---NDU
											8 => "0001011011000000",  ---ADI
											9 => "0000100010100001",  ---ADD
											10 => "0000000000000000", ---ADD
											11 => "0010110110110010", ---NDC
											12 => "1100110101111010", ---BEQ
											13 => "0101100101010110", ---SW
											29 => "0001011011000001", ---ADI
											30 => "0001110110010111", ---ADI
											31 => "0101000110000100", ---SW
											32 => "0100000110000000", ---LW
											33 => "0100001110000001", ---LW
											34 => "1100101001001011", ---BEQ
											35 => "0000000010010000", ---ADD
											36 => "0000011100100010", ---ADD
											37 => "0001001001111111", ---ADI
											38 => "0001111111111011", ---ADI
											46 => "0101010110000010", ---SW
											47 => "0101100110000011", ---SW
											48 => "0001011011111111", ---ADI
											49 => "0101011110000101", ---SW
											50 => "0100111110000100", ---LW
											others => "0000000000000000");
begin
	process(clock,mem_Write,mem_read,Din,A,T)
	begin
		if((mem_Write) = '1') then
			T(to_integer(unsigned(A)))<= Din;
		elsif(mem_read = '1') then
			Dout <= T(to_integer(unsigned(A)));
		end if;
	end process;
end Structure;
